library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity Decoder_5_32 is
    Port ( 
        Dec_Awr: in  STD_LOGIC_VECTOR (4 downto 0);
        Dec_Output : out STD_LOGIC_VECTOR(31 downto 0)
    );
end Decoder_5_32;

architecture Behavioral of Decoder_5_32 is

begin

	Dec_Output <= 	"00000000000000000000000000000001"   when Dec_Awr = "00000" else
					"00000000000000000000000000000010"   when Dec_Awr = "00001" else
					"00000000000000000000000000000100"   when Dec_Awr = "00010" else
					"00000000000000000000000000001000"   when Dec_Awr = "00011" else
					"00000000000000000000000000010000"   when Dec_Awr = "00100" else
					"00000000000000000000000000100000"   when Dec_Awr = "00101" else
					"00000000000000000000000001000000"   when Dec_Awr = "00110" else
					"00000000000000000000000010000000"   when Dec_Awr = "00111" else
					"00000000000000000000000100000000"   when Dec_Awr = "01000" else
					"00000000000000000000001000000000"   when Dec_Awr = "01001" else
					"00000000000000000000010000000000"   when Dec_Awr = "01010" else
					"00000000000000000000100000000000"   when Dec_Awr = "01011" else
					"00000000000000000001000000000000"   when Dec_Awr = "01100" else
					"00000000000000000010000000000000"   when Dec_Awr = "01101" else
					"00000000000000000100000000000000"   when Dec_Awr = "01110" else
					"00000000000000001000000000000000"   when Dec_Awr = "01111" else
					"00000000000000010000000000000000"   when Dec_Awr = "10000" else
					"00000000000000100000000000000000"   when Dec_Awr = "10001" else
					"00000000000001000000000000000000"   when Dec_Awr = "10010" else
					"00000000000010000000000000000000"   when Dec_Awr = "10011" else
					"00000000000100000000000000000000"   when Dec_Awr = "10100" else
					"00000000001000000000000000000000"   when Dec_Awr = "10101" else
					"00000000010000000000000000000000"   when Dec_Awr = "10110" else
					"00000000100000000000000000000000"   when Dec_Awr = "10111" else
					"00000001000000000000000000000000"   when Dec_Awr = "11000" else
					"00000010000000000000000000000000"   when Dec_Awr = "11001" else
					"00000100000000000000000000000000"   when Dec_Awr = "11010" else
					"00001000000000000000000000000000"   when Dec_Awr = "11011" else
					"00010000000000000000000000000000"   when Dec_Awr = "11100" else
					"00100000000000000000000000000000"   when Dec_Awr = "11101" else
					"01000000000000000000000000000000"   when Dec_Awr = "11110" else
					"10000000000000000000000000000000";

end Behavioral;